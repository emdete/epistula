module vmime

fn init() {
}
