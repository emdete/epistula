module gmime

fn init() {
}
