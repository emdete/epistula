module vmime

fn init() {
	eprintln("hi from vmime")
}
